`timescale 1ns / 1ps

module addr_counter(

    );
    
endmodule
